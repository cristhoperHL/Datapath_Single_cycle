module Data_memory(address,write_data,Memwrite,Memread,read_data);

input [31:0] address,write_data;
input Memwrite,Memread;
output [31:0] read_data;





endmodule 