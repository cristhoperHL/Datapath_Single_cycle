module Register_file();


endmodule