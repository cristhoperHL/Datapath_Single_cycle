module Data_memory();

endmodule 